library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_ARITH.all;


entity imem is
    port(
         clk      : in  std_ulogic;
         addr     : in  std_ulogic_vector (6 downto 0);
         data     : out std_ulogic_vector (7 downto 0)
         );
end imem;

architecture BHV of imem is

    type ROM_TYPE is array (0 to 127) of std_ulogic_vector (7 downto 0);

    constant rom_content : ROM_TYPE := (
    "10110000", -- IN r0, xx
    "10110100", -- IN r1, xx
    "10111000", -- IN r2, xx
    "10111100", -- IN r3, xx
    "01000001", -- add r0, r1
	"00000000",	 -- nop
	"00000000",  --  nop
	"11111100",
	"00001110",	
	"10000000",	
	"10111111",
	"00001111",	
	"10000000",	
	"10110100",
	--"11100100",	-- commented these out randomly because total must = 127
	--"11110101",	
	--"10000000",
	--"00100010",	 
	"10001011",	
	"00010010",
	"10001010",	
	"00010011",
	"10001001",	
	"00010100",
	"10001101",	
	"00010101",
	"11100100",	
	"11110101",	
	"00010110",
	"10101101",	
	"00010110",
	"11101101",	
	"00110011",	
	"10010101",	
	"11100000",
	"11111100",	
	"11000011",	
	"11101101",	
	"10010101",	
	"00010101",
	"01110100",	
	"10000000",
	"11111000",	
	"01101100",	
	"10011000",	
	"01010000",
	"00011001",
	"10101011",	
	"00010010",
	"10101010",	
	"00010011",
	"10101001",	
	"00010100",
	"10101111",	
	"00010110",
	"11101111",	
	"00110011",	
	"10010101",	
	"11100000",
	"10001111",	
	"10000010",
	"11110101",	
	"10000011",
	"00010010",	
	"00000001",
	"11001111",
	"11110101",	
	"10000000",
	"00000101",	
	"00010110",
	"10000000",	
	"11010101",
	"00100010",	
	"01111000",	
	"00001000",
	"01111100",	
	"00000000",
	"01111101",	
	"00000000",
	"01111011",	
	"11111111",
	"01111010",	
	"00000000",
	"01111001",	
	"11000000",
	"01111110",	
	"00000000",
	"01111111",
	"00001010",
	"00010010",	
	"00000001",
	"10100110",
	"01111011",
	"00000000",
	"01111010",	
	"00000000",
	"01111001",	
	"00001000",
	"01111101",
	"00001010",
	"00010010",	
	"00000000",
	"00000011",
	"01111011",	
	"00000000",
	"01111010",	
	"00000000",
	"01111001",	
	"00001000",
	"01111101",	
	"00001010",
	"00010010",	
	"00000000",
	"01011101",
	"10000000",	
	"11111110",
	"00100010",
	"00010011",	
	"00010010",	
	"00010001",
	"00010000",
	"00001111",	
	"00001110",	
	"00001101",	
	"00001100",	
	"00001011",	
	"00001010",	
	"01111000",	
	"01111111",
	"11100100",	
	"11110110",	
	"11011000");
begin

p1:    process (clk)
	 variable add_in : integer := 0;
    begin
        if rising_edge(clk) then
					 add_in := conv_integer(unsigned(addr));
                data <= rom_content(add_in);
        end if;
    end process;
end BHV;
